* /home/dilip/eSim-Workspace/Mixed_Signal_Based_Buck_Converter/Mixed_Signal_Based_Buck_Converter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Apr 14 19:44:45 2022

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Vin Net-_Q1-Pad2_ Net-_D1-Pad2_ eSim_NPN		
L1  Net-_D1-Pad2_ Vout 1		
D1  GND Net-_D1-Pad2_ eSim_Diode		
C1  Vout GND 10n		
R1  Vout GND 10k		
v2  Vin GND DC		
U6  Vout plot_v1		
U4  Vin plot_v1		
v1  clk GND pulse		
U3  clk Net-_U1-Pad1_ adc_bridge_1		
U5  Net-_U1-Pad2_ Net-_Q1-Pad2_ dac_bridge_1		
U2  clk plot_v1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ pwm		

.end
